CDLv2�H�\                                                                                                                   				  		                                                               		                                                                                                                                                                                                                                                                                                        	                                  	                                                                                        	                                                                 		        	    	  				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    							      				                      	   	                                                                    	                                 				                                                                                                                                                                                                      	                         		                                                                                                             	                                                                                                                                                                                                                                      	                                           		                                                                                                                                                                                                                                                             	                                           				          	             				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            	  		                                                                                                                                                                                                 				                         	                                           	                                     			                    	                                                                                      	                    	                                                                                                                                                     	                                                                                                                                                                                                                                                                     	                                                                                                                                                                                                                                                                                                                                                  		  	         	            		         	                     		                        									                                          	                                                                              	                                                                                                                                                                                                                                                 	           	                                                                                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             	                                                                                                                                          	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      	            	                                                        	                                                                                            	                  		                                                             		         		          	                                                                                                                                                                                                                                                            			                                                                                          		                   	 	                                                                                             	 		     	    	                                                                                                             			                                                                           			                            			               	   		                                    	                     				                                                                                                                                                                                                                                                                                       			                                                                                                                                             	          	                                                                                                                                                                                                                                                                                      	                                                                                                                                                                                                                                                                                    					        			                                                                                                                                                                                                                                             	                                                			                  				          							          	 					 	      										                                                 		                                                                	                        	       			    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     