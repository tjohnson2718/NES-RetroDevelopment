CDLv2�H�\                                                                                                                   				    		                                                                                                     	          	                                                                                                                                                                                                                                                                                                        	                                         	                                                                                                                                           	                                                                           		            	                            				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    							      				               	     	                                                                                                                                                                 	                                 				                                                                                                                                                                                                                                                                               		                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 	                                                                                                                                                                                                                                                                                                                                                        	                                           			                  	             				                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   			                                                                                                                                                                                                                                                                  	   	                                                                                                                                     	                                                                                                                                        	                                                                          			                                                                                                                                                                                                                                                                                              	                             	                                                                                                                                                       	                                                                                                                                                                                                                                                                                                                                                           	                                                                                                                                                                                                                                                                                                                                                                             	  	         	            			 	  		                    			             						                                    	    	                                                                              	                                                                                                                                                                                                                                         		                                                                                                                                                                                         	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  	                                                                                                                                          	                                                                                                                                                                                                                                    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               	               	                                                             		         		                                                                          	                                                                                                                                                                                                                                                            			                                                                                                                                                                                                                                                             		                   	 	                                                                                             	 		     	     	                                    	                                                                                          				                                         		                                                                                              		               	   		                                                  				                                                                                                                                                                                                                                                                                                                                                                                                   		                                                                                                                                             	     	                                                                                                                                                                                                                                                                                            	                                                                                                                                                                                                                                                                                    					                 			                                                                                                                                                                                                                                                                                                                                                                                                                    	                                                                                     			                                				                 					                    	  					    	      								                    	              	                                                     		                                                                	                        	          			    	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       